library ieee;
use ieee.std_logic_1164.all;

--! \memorymap external example.toml
entity example is
    port (
        clock : in  std_logic;
        reset : in  std_logic
    );
end entity example;
